module adder ( input bit[3:0] a, b, output bit[4:0] c );

	assign c = a + b;

endmodule

